`timescale 1ns / 1ps
`include "include.v"

module Weight_Memory #(
    //numWeight: 
    parameter numWeight = 3, neuronNo = 1, layerNo = 1, addressWidth = 10, dataWidth = 16, weightFile = "w_1_15.mif"
) (
    input clk,
    input wen,
    input ren,
    input [addressWidth-1 : 0] wadd,
    input [addressWidth-1 : 0] radd,
    input [dataWidth-1 : 0] win,
    output reg [dataWidth-1 : 0] wout);

    reg [dataWidth-1 : 0] mem [numWeight-1 : 0];    //numWeight个 位宽为dataWidth的 一维数组

    `ifdef pretrained
        initial
            begin
                $readmemb(weightFile, mem);
            end
        `else
            always @(posedge clk) begin
                if(wen)
                begin
                    mem[wadd] <= win;
                end
            end
    `endif 

    always @(posedge clk) begin
        if (ren) begin
            wout <= mem[radd];
        end
    end
    
endmodule